magic
tech siliwiz
magscale 1 1
timestamp 1750324749
<< pmos >>
rect 8 1 392 384
<< nwell >>
rect 96 223 305 372
rect 95 221 349 377
<< ndiffusion >>
rect 132 85 270 131
<< pdiffusion >>
rect 132 254 270 316
<< psubstratepdiff >>
rect 319 0 382 58
<< nsubstratendiff >>
rect 291 309 338 361
<< polysilicon >>
rect 178 51 217 327
rect 148 179 201 220
<< pdcontact >>
rect 233 264 266 307
rect 132 259 169 312
<< ndcontact >>
rect 236 89 268 127
rect 132 88 166 128
<< polycontact >>
rect 147 185 172 214
<< nsubstratencontact >>
rect 295 330 335 364
<< psubstratepcontact >>
rect 333 8 377 49
<< metal1 >>
rect 39 179 127 218
rect 270 180 366 218
rect 110 179 173 216
rect 229 89 270 307
rect 244 180 284 214
rect 128 264 164 366
rect 132 13 166 130
rect 40 9 374 49
rect 42 334 358 373
rect 29 328 80 377
rect 30 6 81 56
<< labels >>
flabel pmos s 8 1 392 384 0 FreeSans 240 90 0 0 
port 1 nsew signal output
flabel metal1 s 39 179 127 218 0 FreeSans 240 90 0 0 in
port 2 nsew signal output
flabel metal1 s 270 180 366 218 0 FreeSans 240 90 0 0 out
port 3 nsew signal output
flabel metal1 s 29 328 80 377 0 FreeSans 240 90 0 0 vdd
port 4 nsew signal output
flabel metal1 s 30 6 81 56 0 FreeSans 240 90 0 0 vss
port 5 nsew signal output
<< end >>